module nexysVideo (
    input clk
);

endmodule
